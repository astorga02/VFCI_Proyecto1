class Generador#(parameter message, tama_de_paquete,controladores,caso,opcion,broadcast);
  
endclass
